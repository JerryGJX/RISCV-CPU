`include "definition.v"


module insFetcher(
    input wire clk,
    input wire rst,
    input wire rdy,

    
);