
module memCtrl(
    input wire clk,
    input wire rst,
    input wire rdy,

    input wire clr,

    
)