// `ifndef _predictor
// `define _predictor
// `include "definition.v"

// module predictor (
//     input wire clk,
//     input wire rst,
//     input wire rdy,
//     input wire rollback,

//     //with ifetch
//     input  wire                query_enable,
//     input  wire [`OPENUM_TYPE] op_enum,
//     input  wire [  `ADDR_TYPE] now_pc,
//     output reg  [  `ADDR_TYPE] next_pc,
//     output reg                 inst_pred_jump,


//     //with rob
//     input wire rob_br_commit,
//     input wire rob_br_jump
// );

// endmodule
// `endif
