`ifndef macro_rs
`define macro_rs
`include "definition.v"

module RS (
    input wire clk,
    input wire rst,
    input wire rdy,

    //RS
    output reg RS_next_full

);

endmodule
`endif
