`include "riscv/src/definition.v"

module RS(
    input wire clk,
    input wire rst,
    input wire clr,
    input wire rdy,

    //RS
    output reg RS_next_full,
    output reg [`]


);

endmodule